/******************************************************************************
 * (C) Copyright 2015 AMIQ Consulting
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * MODULE:      scrambler_descrambler_types.svh
 * PROJECT:     scrambler_descrambler
 *
 *
 * Description: This is the file with the types used by the package
 *******************************************************************************/


`ifndef SCRAMBLER_DESCRAMBLER_TYPES_SVH
`define SCRAMBLER_DESCRAMBLER_TYPES_SVH


// unpacked array of bits to model streams of bits
typedef bit bs_t[];


`endif