/******************************************************************************
 * (C) Copyright 2015 AMIQ Consulting
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * MODULE:      scrambler_descrambler_pkg.sv
 * PROJECT:     scrambler_descrambler
 *
 *
 * Description: This is the package file
 *******************************************************************************/

`ifndef SCRAMBLER_DESCRAMBLER_PKG_SV
`define SCRAMBLER_DESCRAMBLER_PKG_SV

package scrambler_descrambler_pkg;
   import uvm_pkg::*;
   `include "uvm_macros.svh"

   `include "scrambler_descrambler_types.svh";
   `include "scrambler_descrambler_additive.svh";
   `include "scrambler_multiplicative.svh";
   `include "descrambler_multiplicative.svh";

endpackage

`endif//SCRAMBLER_DESCRAMBLER_PKG_SV